`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer: 
// 
// Create Date: 2021/06/19 21:27:33
// Design Name: 
// Module Name: mul_16x256
// Project Name: 
// Target Devices: 
// Tool Versions: 
// Description: 
// 
// Dependencies: 
// 
// Revision:
// Revision 0.01 - File Created
// Additional Comments:
// 
//////////////////////////////////////////////////////////////////////////////////


module mul_16x256(
    input   wire    clk,
    input   wire    reset,
    input   wire    [15:0]a,
    input   wire    [255:0]b,
    output  reg     [271:0]out,
    output  reg     done
    );
    
    
    
endmodule
