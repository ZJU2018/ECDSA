`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer: 
// 
// Create Date: 2021/04/15 15:01:12
// Design Name: 
// Module Name: hash
// Project Name: 
// Target Devices: 
// Tool Versions: 
// Description: hash the message
// sha-1
// Dependencies: 
// 
// Revision:
// Revision 0.01 - File Created
// Additional Comments:
// 
//////////////////////////////////////////////////////////////////////////////////
module hash(
    input   wire    clk,
    input   wire    reset,
    input   wire    start,
    input   wire    [512:0] in,
    output  wire    [159:0] hash,
    output  reg     done
    );

    reg [31:0]AA, A;
    reg [31:0]BB, B;
    reg [31:0]CC, C;
    reg [31:0]DD, D;
    reg [31:0]EE, E;
    wire [31:0]W[0:79];
    reg [6:0]count;
    
    assign W[0] = in[511:480];
    assign W[1] = in[479:448];
    assign W[2] = in[447:416];
    assign W[3] = in[415:384];
    assign W[4] = in[383:352];
    assign W[5] = in[351:320];
    assign W[6] = in[319:288];
    assign W[7] = in[287:256];
    assign W[8] = in[255:224];
    assign W[9] = in[223:192];
    assign W[10] = in[191:160];
    assign W[11] = in[159:128];
    assign W[12] = in[127:96];
    assign W[13] = in[95:64];
    assign W[14] = in[63:32];
    assign W[15] = in[31:0];
    assign W[16] = {W[13][30:0],W[13][31]} ^ {W[8][30:0],W[8][31]} ^ {W[2][30:0],W[2][31]} ^ {W[0][30:0],W[0][31]};
    assign W[17] = {W[14][30:0],W[14][31]} ^ {W[9][30:0],W[9][31]} ^ {W[3][30:0],W[3][31]} ^ {W[1][30:0],W[1][31]};
    assign W[18] = {W[15][30:0],W[15][31]} ^ {W[10][30:0],W[10][31]} ^ {W[4][30:0],W[4][31]} ^ {W[2][30:0],W[2][31]};
    assign W[19] = {W[16][30:0],W[16][31]} ^ {W[11][30:0],W[11][31]} ^ {W[5][30:0],W[5][31]} ^ {W[3][30:0],W[3][31]};
    assign W[20] = {W[17][30:0],W[17][31]} ^ {W[12][30:0],W[12][31]} ^ {W[6][30:0],W[6][31]} ^ {W[4][30:0],W[4][31]};
    assign W[21] = {W[18][30:0],W[18][31]} ^ {W[13][30:0],W[13][31]} ^ {W[7][30:0],W[7][31]} ^ {W[5][30:0],W[5][31]};
    assign W[22] = {W[19][30:0],W[19][31]} ^ {W[14][30:0],W[14][31]} ^ {W[8][30:0],W[8][31]} ^ {W[6][30:0],W[6][31]};
    assign W[23] = {W[20][30:0],W[20][31]} ^ {W[15][30:0],W[15][31]} ^ {W[9][30:0],W[9][31]} ^ {W[7][30:0],W[7][31]};
    assign W[24] = {W[21][30:0],W[21][31]} ^ {W[16][30:0],W[16][31]} ^ {W[10][30:0],W[10][31]} ^ {W[8][30:0],W[8][31]};
    assign W[25] = {W[22][30:0],W[22][31]} ^ {W[17][30:0],W[17][31]} ^ {W[11][30:0],W[11][31]} ^ {W[9][30:0],W[9][31]};
    assign W[26] = {W[23][30:0],W[23][31]} ^ {W[18][30:0],W[18][31]} ^ {W[12][30:0],W[12][31]} ^ {W[10][30:0],W[10][31]};
    assign W[27] = {W[24][30:0],W[24][31]} ^ {W[19][30:0],W[19][31]} ^ {W[13][30:0],W[13][31]} ^ {W[11][30:0],W[11][31]};
    assign W[28] = {W[25][30:0],W[25][31]} ^ {W[20][30:0],W[20][31]} ^ {W[14][30:0],W[14][31]} ^ {W[12][30:0],W[12][31]};
    assign W[29] = {W[26][30:0],W[26][31]} ^ {W[21][30:0],W[21][31]} ^ {W[15][30:0],W[15][31]} ^ {W[13][30:0],W[13][31]};
    assign W[30] = {W[27][30:0],W[27][31]} ^ {W[22][30:0],W[22][31]} ^ {W[16][30:0],W[16][31]} ^ {W[14][30:0],W[14][31]};
    assign W[31] = {W[28][30:0],W[28][31]} ^ {W[23][30:0],W[23][31]} ^ {W[17][30:0],W[17][31]} ^ {W[15][30:0],W[15][31]};
    assign W[32] = {W[29][30:0],W[29][31]} ^ {W[24][30:0],W[24][31]} ^ {W[18][30:0],W[18][31]} ^ {W[16][30:0],W[16][31]};
    assign W[33] = {W[30][30:0],W[30][31]} ^ {W[25][30:0],W[25][31]} ^ {W[19][30:0],W[19][31]} ^ {W[17][30:0],W[17][31]};
    assign W[34] = {W[31][30:0],W[31][31]} ^ {W[26][30:0],W[26][31]} ^ {W[20][30:0],W[20][31]} ^ {W[18][30:0],W[18][31]};
    assign W[35] = {W[32][30:0],W[32][31]} ^ {W[27][30:0],W[27][31]} ^ {W[21][30:0],W[21][31]} ^ {W[19][30:0],W[19][31]};
    assign W[36] = {W[33][30:0],W[33][31]} ^ {W[28][30:0],W[28][31]} ^ {W[22][30:0],W[22][31]} ^ {W[20][30:0],W[20][31]};
    assign W[37] = {W[34][30:0],W[34][31]} ^ {W[29][30:0],W[29][31]} ^ {W[23][30:0],W[23][31]} ^ {W[21][30:0],W[21][31]};
    assign W[38] = {W[35][30:0],W[35][31]} ^ {W[30][30:0],W[30][31]} ^ {W[24][30:0],W[24][31]} ^ {W[22][30:0],W[22][31]};
    assign W[39] = {W[36][30:0],W[36][31]} ^ {W[31][30:0],W[31][31]} ^ {W[25][30:0],W[25][31]} ^ {W[23][30:0],W[23][31]};
    assign W[40] = {W[37][30:0],W[37][31]} ^ {W[32][30:0],W[32][31]} ^ {W[26][30:0],W[26][31]} ^ {W[24][30:0],W[24][31]};
    assign W[41] = {W[38][30:0],W[38][31]} ^ {W[33][30:0],W[33][31]} ^ {W[27][30:0],W[27][31]} ^ {W[25][30:0],W[25][31]};
    assign W[42] = {W[39][30:0],W[39][31]} ^ {W[34][30:0],W[34][31]} ^ {W[28][30:0],W[28][31]} ^ {W[26][30:0],W[26][31]};
    assign W[43] = {W[40][30:0],W[40][31]} ^ {W[35][30:0],W[35][31]} ^ {W[29][30:0],W[29][31]} ^ {W[27][30:0],W[27][31]};
    assign W[44] = {W[41][30:0],W[41][31]} ^ {W[36][30:0],W[36][31]} ^ {W[30][30:0],W[30][31]} ^ {W[28][30:0],W[28][31]};
    assign W[45] = {W[42][30:0],W[42][31]} ^ {W[37][30:0],W[37][31]} ^ {W[31][30:0],W[31][31]} ^ {W[29][30:0],W[29][31]};
    assign W[46] = {W[43][30:0],W[43][31]} ^ {W[38][30:0],W[38][31]} ^ {W[32][30:0],W[32][31]} ^ {W[30][30:0],W[30][31]};
    assign W[47] = {W[44][30:0],W[44][31]} ^ {W[39][30:0],W[39][31]} ^ {W[33][30:0],W[33][31]} ^ {W[31][30:0],W[31][31]};
    assign W[48] = {W[45][30:0],W[45][31]} ^ {W[40][30:0],W[40][31]} ^ {W[34][30:0],W[34][31]} ^ {W[32][30:0],W[32][31]};
    assign W[49] = {W[46][30:0],W[46][31]} ^ {W[41][30:0],W[41][31]} ^ {W[35][30:0],W[35][31]} ^ {W[33][30:0],W[33][31]};
    assign W[50] = {W[47][30:0],W[47][31]} ^ {W[42][30:0],W[42][31]} ^ {W[36][30:0],W[36][31]} ^ {W[34][30:0],W[34][31]};
    assign W[51] = {W[48][30:0],W[48][31]} ^ {W[43][30:0],W[43][31]} ^ {W[37][30:0],W[37][31]} ^ {W[35][30:0],W[35][31]};
    assign W[52] = {W[49][30:0],W[49][31]} ^ {W[44][30:0],W[44][31]} ^ {W[38][30:0],W[38][31]} ^ {W[36][30:0],W[36][31]};
    assign W[53] = {W[50][30:0],W[50][31]} ^ {W[45][30:0],W[45][31]} ^ {W[39][30:0],W[39][31]} ^ {W[37][30:0],W[37][31]};
    assign W[54] = {W[51][30:0],W[51][31]} ^ {W[46][30:0],W[46][31]} ^ {W[40][30:0],W[40][31]} ^ {W[38][30:0],W[38][31]};
    assign W[55] = {W[52][30:0],W[52][31]} ^ {W[47][30:0],W[47][31]} ^ {W[41][30:0],W[41][31]} ^ {W[39][30:0],W[39][31]};
    assign W[56] = {W[53][30:0],W[53][31]} ^ {W[48][30:0],W[48][31]} ^ {W[42][30:0],W[42][31]} ^ {W[40][30:0],W[40][31]};
    assign W[57] = {W[54][30:0],W[54][31]} ^ {W[49][30:0],W[49][31]} ^ {W[43][30:0],W[43][31]} ^ {W[41][30:0],W[41][31]};
    assign W[58] = {W[55][30:0],W[55][31]} ^ {W[50][30:0],W[50][31]} ^ {W[44][30:0],W[44][31]} ^ {W[42][30:0],W[42][31]};
    assign W[59] = {W[56][30:0],W[56][31]} ^ {W[51][30:0],W[51][31]} ^ {W[45][30:0],W[45][31]} ^ {W[43][30:0],W[43][31]};
    assign W[60] = {W[57][30:0],W[57][31]} ^ {W[52][30:0],W[52][31]} ^ {W[46][30:0],W[46][31]} ^ {W[44][30:0],W[44][31]};
    assign W[61] = {W[58][30:0],W[58][31]} ^ {W[53][30:0],W[53][31]} ^ {W[47][30:0],W[47][31]} ^ {W[45][30:0],W[45][31]};
    assign W[62] = {W[59][30:0],W[59][31]} ^ {W[54][30:0],W[54][31]} ^ {W[48][30:0],W[48][31]} ^ {W[46][30:0],W[46][31]};
    assign W[63] = {W[60][30:0],W[60][31]} ^ {W[55][30:0],W[55][31]} ^ {W[49][30:0],W[49][31]} ^ {W[47][30:0],W[47][31]};
    assign W[64] = {W[61][30:0],W[61][31]} ^ {W[56][30:0],W[56][31]} ^ {W[50][30:0],W[50][31]} ^ {W[48][30:0],W[48][31]};
    assign W[65] = {W[62][30:0],W[62][31]} ^ {W[57][30:0],W[57][31]} ^ {W[51][30:0],W[51][31]} ^ {W[49][30:0],W[49][31]};
    assign W[66] = {W[63][30:0],W[63][31]} ^ {W[58][30:0],W[58][31]} ^ {W[52][30:0],W[52][31]} ^ {W[50][30:0],W[50][31]};
    assign W[67] = {W[64][30:0],W[64][31]} ^ {W[59][30:0],W[59][31]} ^ {W[53][30:0],W[53][31]} ^ {W[51][30:0],W[51][31]};
    assign W[68] = {W[65][30:0],W[65][31]} ^ {W[60][30:0],W[60][31]} ^ {W[54][30:0],W[54][31]} ^ {W[52][30:0],W[52][31]};
    assign W[69] = {W[66][30:0],W[66][31]} ^ {W[61][30:0],W[61][31]} ^ {W[55][30:0],W[55][31]} ^ {W[53][30:0],W[53][31]};
    assign W[70] = {W[67][30:0],W[67][31]} ^ {W[62][30:0],W[62][31]} ^ {W[56][30:0],W[56][31]} ^ {W[54][30:0],W[54][31]};
    assign W[71] = {W[68][30:0],W[68][31]} ^ {W[63][30:0],W[63][31]} ^ {W[57][30:0],W[57][31]} ^ {W[55][30:0],W[55][31]};
    assign W[72] = {W[69][30:0],W[69][31]} ^ {W[64][30:0],W[64][31]} ^ {W[58][30:0],W[58][31]} ^ {W[56][30:0],W[56][31]};
    assign W[73] = {W[70][30:0],W[70][31]} ^ {W[65][30:0],W[65][31]} ^ {W[59][30:0],W[59][31]} ^ {W[57][30:0],W[57][31]};
    assign W[74] = {W[71][30:0],W[71][31]} ^ {W[66][30:0],W[66][31]} ^ {W[60][30:0],W[60][31]} ^ {W[58][30:0],W[58][31]};
    assign W[75] = {W[72][30:0],W[72][31]} ^ {W[67][30:0],W[67][31]} ^ {W[61][30:0],W[61][31]} ^ {W[59][30:0],W[59][31]};
    assign W[76] = {W[73][30:0],W[73][31]} ^ {W[68][30:0],W[68][31]} ^ {W[62][30:0],W[62][31]} ^ {W[60][30:0],W[60][31]};
    assign W[77] = {W[74][30:0],W[74][31]} ^ {W[69][30:0],W[69][31]} ^ {W[63][30:0],W[63][31]} ^ {W[61][30:0],W[61][31]};
    assign W[78] = {W[75][30:0],W[75][31]} ^ {W[70][30:0],W[70][31]} ^ {W[64][30:0],W[64][31]} ^ {W[62][30:0],W[62][31]};
    assign W[79] = {W[76][30:0],W[76][31]} ^ {W[71][30:0],W[71][31]} ^ {W[65][30:0],W[65][31]} ^ {W[63][30:0],W[63][31]};
    assign hash = {A,B,C,D,E};
    
    always@(posedge clk or negedge reset)begin
        if(~reset)begin
            A <= 32'h67452301;
            B <= 32'hEFCDAB89;
            C <= 32'h98BADCFE;
            D <= 32'h10325476;
            E <= 32'hC3D2E1F0;
        end
        else if(start)begin
            A <= A;
            B <= B;
            C <= C;
            D <= D;
            E <= E;
        end 
        else begin
            if(count < 20)begin
                A <= {A[26:0],A[31:27]} + ((B & C) | (~B & D)) + E + W[count] + 32'h5A827999;
                B <= A;
                C <= {B[1:0],B[31:2]};
                D <= C;
                E <= D;
            end
            else if(count < 40)begin
                A <= {A[26:0],A[31:27]} + (B ^ C ^ D) + E + W[count] + 32'h6ED9EBA1;
                B <= A;
                C <= {B[1:0],B[31:2]};
                D <= C;
                E <= D;
            end
            else if(count < 60)begin
                A <= {A[26:0],A[31:27]} + ((B & C) | (B & D) | (C & D)) + E + W[count] + 32'h8F1BBCDC;
                B <= A;
                C <= {B[1:0],B[31:2]};
                D <= C;
                E <= D;
            end
            else if(count < 80)begin
                A <= {A[26:0],A[31:27]} + (B ^ C ^ D) + E + W[count] + 32'hCA62C1D6;
                B <= A;
                C <= {B[1:0],B[31:2]};
                D <= C;
                E <= D;
            end
            else if(count ==80)begin
                A <= A + AA;
                B <= B + BB;
                C <= C + CC;
                D <= D + DD;
                E <= E + EE;
            end
            else begin
                A <= A;
                B <= B;
                C <= C;
                D <= D;
                E <= E;
            end
        end
    end
    
    
        always@(posedge clk or negedge reset)begin
        if(~reset)begin
            AA <= 32'h67452301;
            BB <= 32'hEFCDAB89;
            CC <= 32'h98BADCFE;
            DD <= 32'h10325476;
            EE <= 32'hC3D2E1F0;
        end
        else if(done)begin
            AA <= A;
            BB <= B;
            CC <= C;
            DD <= D;
            EE <= E;
        end
    end

    always@(posedge clk or negedge reset)begin
        if(~reset)begin
            count <= 0;
        end
        else if(start)begin
            count <= 0;
        end
        else if(count <=80)begin
            count <= count + 1;
        end
        else
            count <= count;  
    end
    
    always@(posedge clk or negedge reset)begin
        if(~reset)begin
            done <= 0;
        end 
        else if(count == 80)begin
            done <= 1;
        end
        else begin
            done <= 0;
        end
    end
    
endmodule
